module conv2d_4(                               
     input wire clk,                                             
     input wire rst,                                             
     input wire load,                                             
     input wire input_valid,                                             
     input wire sof,                                             
     output wire o_sof,                                             
     output wire load_success,                                             
     output wire output_valid,                                      
     output wire [31:0] d_out[15:0],    
     input wire [31:0] d_in[7:0]                    
); 
wire output_valid_affter_conv;                                             
wire [31:0] _0_addbus_[7:0];    
conv2d #("weight/conv2d_4/0_0.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_0_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(load_success),
	.output_valid(output_valid_affter_conv),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_0_addbus_[0])
);
conv2d #("weight/conv2d_4/0_1.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_0_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_0_addbus_[1])
);
conv2d #("weight/conv2d_4/0_2.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_0_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_0_addbus_[2])
);
conv2d #("weight/conv2d_4/0_3.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_0_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_0_addbus_[3])
);
conv2d #("weight/conv2d_4/0_4.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_0_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_0_addbus_[4])
);
conv2d #("weight/conv2d_4/0_5.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_0_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_0_addbus_[5])
);
conv2d #("weight/conv2d_4/0_6.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_0_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_0_addbus_[6])
);
conv2d #("weight/conv2d_4/0_7.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_0_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_0_addbus_[7])
);
sum_8 #(3) sum_0( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .output_valid(output_valid), 
        .o_sof(o_sof), 
        .data_out(d_out[0]), 
        .data_in_0(_0_addbus_[0]), 
        .data_in_1(_0_addbus_[1]), 
        .data_in_2(_0_addbus_[2]), 
        .data_in_3(_0_addbus_[3]), 
        .data_in_4(_0_addbus_[4]), 
        .data_in_5(_0_addbus_[5]), 
        .data_in_6(_0_addbus_[6]), 
        .data_in_7(_0_addbus_[7]) 
); 
wire [31:0] _1_addbus_[7:0];    
conv2d #("weight/conv2d_4/1_0.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_1_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_1_addbus_[0])
);
conv2d #("weight/conv2d_4/1_1.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_1_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_1_addbus_[1])
);
conv2d #("weight/conv2d_4/1_2.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_1_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_1_addbus_[2])
);
conv2d #("weight/conv2d_4/1_3.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_1_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_1_addbus_[3])
);
conv2d #("weight/conv2d_4/1_4.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_1_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_1_addbus_[4])
);
conv2d #("weight/conv2d_4/1_5.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_1_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_1_addbus_[5])
);
conv2d #("weight/conv2d_4/1_6.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_1_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_1_addbus_[6])
);
conv2d #("weight/conv2d_4/1_7.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_1_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_1_addbus_[7])
);
sum_8 #(3) sum_1( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[1]), 
        .data_in_0(_1_addbus_[0]), 
        .data_in_1(_1_addbus_[1]), 
        .data_in_2(_1_addbus_[2]), 
        .data_in_3(_1_addbus_[3]), 
        .data_in_4(_1_addbus_[4]), 
        .data_in_5(_1_addbus_[5]), 
        .data_in_6(_1_addbus_[6]), 
        .data_in_7(_1_addbus_[7]) 
); 
wire [31:0] _2_addbus_[7:0];    
conv2d #("weight/conv2d_4/2_0.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_2_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_2_addbus_[0])
);
conv2d #("weight/conv2d_4/2_1.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_2_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_2_addbus_[1])
);
conv2d #("weight/conv2d_4/2_2.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_2_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_2_addbus_[2])
);
conv2d #("weight/conv2d_4/2_3.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_2_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_2_addbus_[3])
);
conv2d #("weight/conv2d_4/2_4.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_2_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_2_addbus_[4])
);
conv2d #("weight/conv2d_4/2_5.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_2_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_2_addbus_[5])
);
conv2d #("weight/conv2d_4/2_6.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_2_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_2_addbus_[6])
);
conv2d #("weight/conv2d_4/2_7.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_2_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_2_addbus_[7])
);
sum_8 #(3) sum_2( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[2]), 
        .data_in_0(_2_addbus_[0]), 
        .data_in_1(_2_addbus_[1]), 
        .data_in_2(_2_addbus_[2]), 
        .data_in_3(_2_addbus_[3]), 
        .data_in_4(_2_addbus_[4]), 
        .data_in_5(_2_addbus_[5]), 
        .data_in_6(_2_addbus_[6]), 
        .data_in_7(_2_addbus_[7]) 
); 
wire [31:0] _3_addbus_[7:0];    
conv2d #("weight/conv2d_4/3_0.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_3_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_3_addbus_[0])
);
conv2d #("weight/conv2d_4/3_1.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_3_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_3_addbus_[1])
);
conv2d #("weight/conv2d_4/3_2.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_3_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_3_addbus_[2])
);
conv2d #("weight/conv2d_4/3_3.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_3_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_3_addbus_[3])
);
conv2d #("weight/conv2d_4/3_4.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_3_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_3_addbus_[4])
);
conv2d #("weight/conv2d_4/3_5.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_3_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_3_addbus_[5])
);
conv2d #("weight/conv2d_4/3_6.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_3_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_3_addbus_[6])
);
conv2d #("weight/conv2d_4/3_7.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_3_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_3_addbus_[7])
);
sum_8 #(3) sum_3( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[3]), 
        .data_in_0(_3_addbus_[0]), 
        .data_in_1(_3_addbus_[1]), 
        .data_in_2(_3_addbus_[2]), 
        .data_in_3(_3_addbus_[3]), 
        .data_in_4(_3_addbus_[4]), 
        .data_in_5(_3_addbus_[5]), 
        .data_in_6(_3_addbus_[6]), 
        .data_in_7(_3_addbus_[7]) 
); 
wire [31:0] _4_addbus_[7:0];    
conv2d #("weight/conv2d_4/4_0.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_4_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_4_addbus_[0])
);
conv2d #("weight/conv2d_4/4_1.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_4_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_4_addbus_[1])
);
conv2d #("weight/conv2d_4/4_2.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_4_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_4_addbus_[2])
);
conv2d #("weight/conv2d_4/4_3.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_4_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_4_addbus_[3])
);
conv2d #("weight/conv2d_4/4_4.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_4_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_4_addbus_[4])
);
conv2d #("weight/conv2d_4/4_5.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_4_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_4_addbus_[5])
);
conv2d #("weight/conv2d_4/4_6.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_4_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_4_addbus_[6])
);
conv2d #("weight/conv2d_4/4_7.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_4_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_4_addbus_[7])
);
sum_8 #(3) sum_4( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[4]), 
        .data_in_0(_4_addbus_[0]), 
        .data_in_1(_4_addbus_[1]), 
        .data_in_2(_4_addbus_[2]), 
        .data_in_3(_4_addbus_[3]), 
        .data_in_4(_4_addbus_[4]), 
        .data_in_5(_4_addbus_[5]), 
        .data_in_6(_4_addbus_[6]), 
        .data_in_7(_4_addbus_[7]) 
); 
wire [31:0] _5_addbus_[7:0];    
conv2d #("weight/conv2d_4/5_0.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_5_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_5_addbus_[0])
);
conv2d #("weight/conv2d_4/5_1.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_5_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_5_addbus_[1])
);
conv2d #("weight/conv2d_4/5_2.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_5_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_5_addbus_[2])
);
conv2d #("weight/conv2d_4/5_3.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_5_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_5_addbus_[3])
);
conv2d #("weight/conv2d_4/5_4.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_5_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_5_addbus_[4])
);
conv2d #("weight/conv2d_4/5_5.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_5_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_5_addbus_[5])
);
conv2d #("weight/conv2d_4/5_6.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_5_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_5_addbus_[6])
);
conv2d #("weight/conv2d_4/5_7.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_5_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_5_addbus_[7])
);
sum_8 #(3) sum_5( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[5]), 
        .data_in_0(_5_addbus_[0]), 
        .data_in_1(_5_addbus_[1]), 
        .data_in_2(_5_addbus_[2]), 
        .data_in_3(_5_addbus_[3]), 
        .data_in_4(_5_addbus_[4]), 
        .data_in_5(_5_addbus_[5]), 
        .data_in_6(_5_addbus_[6]), 
        .data_in_7(_5_addbus_[7]) 
); 
wire [31:0] _6_addbus_[7:0];    
conv2d #("weight/conv2d_4/6_0.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_6_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_6_addbus_[0])
);
conv2d #("weight/conv2d_4/6_1.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_6_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_6_addbus_[1])
);
conv2d #("weight/conv2d_4/6_2.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_6_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_6_addbus_[2])
);
conv2d #("weight/conv2d_4/6_3.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_6_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_6_addbus_[3])
);
conv2d #("weight/conv2d_4/6_4.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_6_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_6_addbus_[4])
);
conv2d #("weight/conv2d_4/6_5.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_6_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_6_addbus_[5])
);
conv2d #("weight/conv2d_4/6_6.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_6_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_6_addbus_[6])
);
conv2d #("weight/conv2d_4/6_7.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_6_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_6_addbus_[7])
);
sum_8 #(3) sum_6( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[6]), 
        .data_in_0(_6_addbus_[0]), 
        .data_in_1(_6_addbus_[1]), 
        .data_in_2(_6_addbus_[2]), 
        .data_in_3(_6_addbus_[3]), 
        .data_in_4(_6_addbus_[4]), 
        .data_in_5(_6_addbus_[5]), 
        .data_in_6(_6_addbus_[6]), 
        .data_in_7(_6_addbus_[7]) 
); 
wire [31:0] _7_addbus_[7:0];    
conv2d #("weight/conv2d_4/7_0.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_7_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_7_addbus_[0])
);
conv2d #("weight/conv2d_4/7_1.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_7_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_7_addbus_[1])
);
conv2d #("weight/conv2d_4/7_2.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_7_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_7_addbus_[2])
);
conv2d #("weight/conv2d_4/7_3.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_7_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_7_addbus_[3])
);
conv2d #("weight/conv2d_4/7_4.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_7_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_7_addbus_[4])
);
conv2d #("weight/conv2d_4/7_5.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_7_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_7_addbus_[5])
);
conv2d #("weight/conv2d_4/7_6.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_7_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_7_addbus_[6])
);
conv2d #("weight/conv2d_4/7_7.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_7_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_7_addbus_[7])
);
sum_8 #(3) sum_7( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[7]), 
        .data_in_0(_7_addbus_[0]), 
        .data_in_1(_7_addbus_[1]), 
        .data_in_2(_7_addbus_[2]), 
        .data_in_3(_7_addbus_[3]), 
        .data_in_4(_7_addbus_[4]), 
        .data_in_5(_7_addbus_[5]), 
        .data_in_6(_7_addbus_[6]), 
        .data_in_7(_7_addbus_[7]) 
); 
wire [31:0] _8_addbus_[7:0];    
conv2d #("weight/conv2d_4/8_0.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_8_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_8_addbus_[0])
);
conv2d #("weight/conv2d_4/8_1.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_8_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_8_addbus_[1])
);
conv2d #("weight/conv2d_4/8_2.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_8_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_8_addbus_[2])
);
conv2d #("weight/conv2d_4/8_3.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_8_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_8_addbus_[3])
);
conv2d #("weight/conv2d_4/8_4.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_8_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_8_addbus_[4])
);
conv2d #("weight/conv2d_4/8_5.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_8_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_8_addbus_[5])
);
conv2d #("weight/conv2d_4/8_6.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_8_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_8_addbus_[6])
);
conv2d #("weight/conv2d_4/8_7.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_8_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_8_addbus_[7])
);
sum_8 #(3) sum_8( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[8]), 
        .data_in_0(_8_addbus_[0]), 
        .data_in_1(_8_addbus_[1]), 
        .data_in_2(_8_addbus_[2]), 
        .data_in_3(_8_addbus_[3]), 
        .data_in_4(_8_addbus_[4]), 
        .data_in_5(_8_addbus_[5]), 
        .data_in_6(_8_addbus_[6]), 
        .data_in_7(_8_addbus_[7]) 
); 
wire [31:0] _9_addbus_[7:0];    
conv2d #("weight/conv2d_4/9_0.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_9_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_9_addbus_[0])
);
conv2d #("weight/conv2d_4/9_1.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_9_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_9_addbus_[1])
);
conv2d #("weight/conv2d_4/9_2.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_9_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_9_addbus_[2])
);
conv2d #("weight/conv2d_4/9_3.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_9_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_9_addbus_[3])
);
conv2d #("weight/conv2d_4/9_4.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_9_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_9_addbus_[4])
);
conv2d #("weight/conv2d_4/9_5.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_9_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_9_addbus_[5])
);
conv2d #("weight/conv2d_4/9_6.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_9_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_9_addbus_[6])
);
conv2d #("weight/conv2d_4/9_7.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_9_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_9_addbus_[7])
);
sum_8 #(3) sum_9( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[9]), 
        .data_in_0(_9_addbus_[0]), 
        .data_in_1(_9_addbus_[1]), 
        .data_in_2(_9_addbus_[2]), 
        .data_in_3(_9_addbus_[3]), 
        .data_in_4(_9_addbus_[4]), 
        .data_in_5(_9_addbus_[5]), 
        .data_in_6(_9_addbus_[6]), 
        .data_in_7(_9_addbus_[7]) 
); 
wire [31:0] _10_addbus_[7:0];    
conv2d #("weight/conv2d_4/10_0.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_10_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_10_addbus_[0])
);
conv2d #("weight/conv2d_4/10_1.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_10_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_10_addbus_[1])
);
conv2d #("weight/conv2d_4/10_2.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_10_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_10_addbus_[2])
);
conv2d #("weight/conv2d_4/10_3.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_10_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_10_addbus_[3])
);
conv2d #("weight/conv2d_4/10_4.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_10_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_10_addbus_[4])
);
conv2d #("weight/conv2d_4/10_5.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_10_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_10_addbus_[5])
);
conv2d #("weight/conv2d_4/10_6.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_10_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_10_addbus_[6])
);
conv2d #("weight/conv2d_4/10_7.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_10_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_10_addbus_[7])
);
sum_8 #(3) sum_10( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[10]), 
        .data_in_0(_10_addbus_[0]), 
        .data_in_1(_10_addbus_[1]), 
        .data_in_2(_10_addbus_[2]), 
        .data_in_3(_10_addbus_[3]), 
        .data_in_4(_10_addbus_[4]), 
        .data_in_5(_10_addbus_[5]), 
        .data_in_6(_10_addbus_[6]), 
        .data_in_7(_10_addbus_[7]) 
); 
wire [31:0] _11_addbus_[7:0];    
conv2d #("weight/conv2d_4/11_0.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_11_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_11_addbus_[0])
);
conv2d #("weight/conv2d_4/11_1.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_11_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_11_addbus_[1])
);
conv2d #("weight/conv2d_4/11_2.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_11_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_11_addbus_[2])
);
conv2d #("weight/conv2d_4/11_3.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_11_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_11_addbus_[3])
);
conv2d #("weight/conv2d_4/11_4.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_11_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_11_addbus_[4])
);
conv2d #("weight/conv2d_4/11_5.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_11_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_11_addbus_[5])
);
conv2d #("weight/conv2d_4/11_6.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_11_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_11_addbus_[6])
);
conv2d #("weight/conv2d_4/11_7.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_11_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_11_addbus_[7])
);
sum_8 #(3) sum_11( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[11]), 
        .data_in_0(_11_addbus_[0]), 
        .data_in_1(_11_addbus_[1]), 
        .data_in_2(_11_addbus_[2]), 
        .data_in_3(_11_addbus_[3]), 
        .data_in_4(_11_addbus_[4]), 
        .data_in_5(_11_addbus_[5]), 
        .data_in_6(_11_addbus_[6]), 
        .data_in_7(_11_addbus_[7]) 
); 
wire [31:0] _12_addbus_[7:0];    
conv2d #("weight/conv2d_4/12_0.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_12_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_12_addbus_[0])
);
conv2d #("weight/conv2d_4/12_1.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_12_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_12_addbus_[1])
);
conv2d #("weight/conv2d_4/12_2.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_12_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_12_addbus_[2])
);
conv2d #("weight/conv2d_4/12_3.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_12_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_12_addbus_[3])
);
conv2d #("weight/conv2d_4/12_4.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_12_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_12_addbus_[4])
);
conv2d #("weight/conv2d_4/12_5.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_12_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_12_addbus_[5])
);
conv2d #("weight/conv2d_4/12_6.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_12_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_12_addbus_[6])
);
conv2d #("weight/conv2d_4/12_7.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_12_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_12_addbus_[7])
);
sum_8 #(3) sum_12( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[12]), 
        .data_in_0(_12_addbus_[0]), 
        .data_in_1(_12_addbus_[1]), 
        .data_in_2(_12_addbus_[2]), 
        .data_in_3(_12_addbus_[3]), 
        .data_in_4(_12_addbus_[4]), 
        .data_in_5(_12_addbus_[5]), 
        .data_in_6(_12_addbus_[6]), 
        .data_in_7(_12_addbus_[7]) 
); 
wire [31:0] _13_addbus_[7:0];    
conv2d #("weight/conv2d_4/13_0.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_13_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_13_addbus_[0])
);
conv2d #("weight/conv2d_4/13_1.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_13_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_13_addbus_[1])
);
conv2d #("weight/conv2d_4/13_2.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_13_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_13_addbus_[2])
);
conv2d #("weight/conv2d_4/13_3.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_13_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_13_addbus_[3])
);
conv2d #("weight/conv2d_4/13_4.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_13_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_13_addbus_[4])
);
conv2d #("weight/conv2d_4/13_5.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_13_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_13_addbus_[5])
);
conv2d #("weight/conv2d_4/13_6.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_13_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_13_addbus_[6])
);
conv2d #("weight/conv2d_4/13_7.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_13_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_13_addbus_[7])
);
sum_8 #(3) sum_13( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[13]), 
        .data_in_0(_13_addbus_[0]), 
        .data_in_1(_13_addbus_[1]), 
        .data_in_2(_13_addbus_[2]), 
        .data_in_3(_13_addbus_[3]), 
        .data_in_4(_13_addbus_[4]), 
        .data_in_5(_13_addbus_[5]), 
        .data_in_6(_13_addbus_[6]), 
        .data_in_7(_13_addbus_[7]) 
); 
wire [31:0] _14_addbus_[7:0];    
conv2d #("weight/conv2d_4/14_0.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_14_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_14_addbus_[0])
);
conv2d #("weight/conv2d_4/14_1.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_14_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_14_addbus_[1])
);
conv2d #("weight/conv2d_4/14_2.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_14_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_14_addbus_[2])
);
conv2d #("weight/conv2d_4/14_3.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_14_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_14_addbus_[3])
);
conv2d #("weight/conv2d_4/14_4.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_14_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_14_addbus_[4])
);
conv2d #("weight/conv2d_4/14_5.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_14_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_14_addbus_[5])
);
conv2d #("weight/conv2d_4/14_6.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_14_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_14_addbus_[6])
);
conv2d #("weight/conv2d_4/14_7.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_14_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_14_addbus_[7])
);
sum_8 #(3) sum_14( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[14]), 
        .data_in_0(_14_addbus_[0]), 
        .data_in_1(_14_addbus_[1]), 
        .data_in_2(_14_addbus_[2]), 
        .data_in_3(_14_addbus_[3]), 
        .data_in_4(_14_addbus_[4]), 
        .data_in_5(_14_addbus_[5]), 
        .data_in_6(_14_addbus_[6]), 
        .data_in_7(_14_addbus_[7]) 
); 
wire [31:0] _15_addbus_[7:0];    
conv2d #("weight/conv2d_4/15_0.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_15_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_15_addbus_[0])
);
conv2d #("weight/conv2d_4/15_1.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_15_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_15_addbus_[1])
);
conv2d #("weight/conv2d_4/15_2.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_15_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_15_addbus_[2])
);
conv2d #("weight/conv2d_4/15_3.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_15_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_15_addbus_[3])
);
conv2d #("weight/conv2d_4/15_4.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_15_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_15_addbus_[4])
);
conv2d #("weight/conv2d_4/15_5.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_15_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_15_addbus_[5])
);
conv2d #("weight/conv2d_4/15_6.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_15_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_15_addbus_[6])
);
conv2d #("weight/conv2d_4/15_7.txt", 0 /*dont use relu*/, 2, 0, 7, 7) conv2d_15_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_15_addbus_[7])
);
sum_8 #(3) sum_15( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[15]), 
        .data_in_0(_15_addbus_[0]), 
        .data_in_1(_15_addbus_[1]), 
        .data_in_2(_15_addbus_[2]), 
        .data_in_3(_15_addbus_[3]), 
        .data_in_4(_15_addbus_[4]), 
        .data_in_5(_15_addbus_[5]), 
        .data_in_6(_15_addbus_[6]), 
        .data_in_7(_15_addbus_[7]) 
); 
endmodule