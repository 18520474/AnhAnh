module conv2d_5(                               
     input wire clk,                                             
     input wire rst,                                             
     input wire load,                                             
     input wire input_valid,                                             
     input wire sof,                                             
     output wire o_sof,                                             
     output wire load_success,                                             
     output wire output_valid,                                      
     output wire [31:0] d_out[15:0],    
     input wire [31:0] d_in[15:0]                    
); 
wire output_valid_affter_conv;                                             
wire [31:0] _0_addbus_[15:0];    
conv2d #("weight/conv2d_5/0_0.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_0_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(load_success),
	.output_valid(output_valid_affter_conv),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_0_addbus_[0])
);
conv2d #("weight/conv2d_5/0_1.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_0_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_0_addbus_[1])
);
conv2d #("weight/conv2d_5/0_2.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_0_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_0_addbus_[2])
);
conv2d #("weight/conv2d_5/0_3.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_0_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_0_addbus_[3])
);
conv2d #("weight/conv2d_5/0_4.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_0_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_0_addbus_[4])
);
conv2d #("weight/conv2d_5/0_5.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_0_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_0_addbus_[5])
);
conv2d #("weight/conv2d_5/0_6.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_0_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_0_addbus_[6])
);
conv2d #("weight/conv2d_5/0_7.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_0_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_0_addbus_[7])
);
conv2d #("weight/conv2d_5/0_8.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_0_8(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[8]),
	.d_out(_0_addbus_[8])
);
conv2d #("weight/conv2d_5/0_9.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_0_9(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[9]),
	.d_out(_0_addbus_[9])
);
conv2d #("weight/conv2d_5/0_10.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_0_10(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[10]),
	.d_out(_0_addbus_[10])
);
conv2d #("weight/conv2d_5/0_11.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_0_11(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[11]),
	.d_out(_0_addbus_[11])
);
conv2d #("weight/conv2d_5/0_12.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_0_12(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[12]),
	.d_out(_0_addbus_[12])
);
conv2d #("weight/conv2d_5/0_13.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_0_13(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[13]),
	.d_out(_0_addbus_[13])
);
conv2d #("weight/conv2d_5/0_14.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_0_14(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[14]),
	.d_out(_0_addbus_[14])
);
conv2d #("weight/conv2d_5/0_15.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_0_15(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[15]),
	.d_out(_0_addbus_[15])
);
sum_16 #(3) sum_0( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .output_valid(output_valid), 
        .o_sof(o_sof), 
        .data_out(d_out[0]), 
        .data_in_0(_0_addbus_[0]), 
        .data_in_1(_0_addbus_[1]), 
        .data_in_2(_0_addbus_[2]), 
        .data_in_3(_0_addbus_[3]), 
        .data_in_4(_0_addbus_[4]), 
        .data_in_5(_0_addbus_[5]), 
        .data_in_6(_0_addbus_[6]), 
        .data_in_7(_0_addbus_[7]), 
        .data_in_8(_0_addbus_[8]), 
        .data_in_9(_0_addbus_[9]), 
        .data_in_10(_0_addbus_[10]), 
        .data_in_11(_0_addbus_[11]), 
        .data_in_12(_0_addbus_[12]), 
        .data_in_13(_0_addbus_[13]), 
        .data_in_14(_0_addbus_[14]), 
        .data_in_15(_0_addbus_[15]) 
); 
wire [31:0] _1_addbus_[15:0];    
conv2d #("weight/conv2d_5/1_0.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_1_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_1_addbus_[0])
);
conv2d #("weight/conv2d_5/1_1.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_1_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_1_addbus_[1])
);
conv2d #("weight/conv2d_5/1_2.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_1_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_1_addbus_[2])
);
conv2d #("weight/conv2d_5/1_3.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_1_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_1_addbus_[3])
);
conv2d #("weight/conv2d_5/1_4.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_1_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_1_addbus_[4])
);
conv2d #("weight/conv2d_5/1_5.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_1_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_1_addbus_[5])
);
conv2d #("weight/conv2d_5/1_6.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_1_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_1_addbus_[6])
);
conv2d #("weight/conv2d_5/1_7.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_1_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_1_addbus_[7])
);
conv2d #("weight/conv2d_5/1_8.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_1_8(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[8]),
	.d_out(_1_addbus_[8])
);
conv2d #("weight/conv2d_5/1_9.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_1_9(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[9]),
	.d_out(_1_addbus_[9])
);
conv2d #("weight/conv2d_5/1_10.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_1_10(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[10]),
	.d_out(_1_addbus_[10])
);
conv2d #("weight/conv2d_5/1_11.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_1_11(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[11]),
	.d_out(_1_addbus_[11])
);
conv2d #("weight/conv2d_5/1_12.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_1_12(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[12]),
	.d_out(_1_addbus_[12])
);
conv2d #("weight/conv2d_5/1_13.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_1_13(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[13]),
	.d_out(_1_addbus_[13])
);
conv2d #("weight/conv2d_5/1_14.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_1_14(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[14]),
	.d_out(_1_addbus_[14])
);
conv2d #("weight/conv2d_5/1_15.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_1_15(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[15]),
	.d_out(_1_addbus_[15])
);
sum_16 #(3) sum_1( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[1]), 
        .data_in_0(_1_addbus_[0]), 
        .data_in_1(_1_addbus_[1]), 
        .data_in_2(_1_addbus_[2]), 
        .data_in_3(_1_addbus_[3]), 
        .data_in_4(_1_addbus_[4]), 
        .data_in_5(_1_addbus_[5]), 
        .data_in_6(_1_addbus_[6]), 
        .data_in_7(_1_addbus_[7]), 
        .data_in_8(_1_addbus_[8]), 
        .data_in_9(_1_addbus_[9]), 
        .data_in_10(_1_addbus_[10]), 
        .data_in_11(_1_addbus_[11]), 
        .data_in_12(_1_addbus_[12]), 
        .data_in_13(_1_addbus_[13]), 
        .data_in_14(_1_addbus_[14]), 
        .data_in_15(_1_addbus_[15]) 
); 
wire [31:0] _2_addbus_[15:0];    
conv2d #("weight/conv2d_5/2_0.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_2_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_2_addbus_[0])
);
conv2d #("weight/conv2d_5/2_1.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_2_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_2_addbus_[1])
);
conv2d #("weight/conv2d_5/2_2.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_2_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_2_addbus_[2])
);
conv2d #("weight/conv2d_5/2_3.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_2_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_2_addbus_[3])
);
conv2d #("weight/conv2d_5/2_4.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_2_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_2_addbus_[4])
);
conv2d #("weight/conv2d_5/2_5.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_2_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_2_addbus_[5])
);
conv2d #("weight/conv2d_5/2_6.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_2_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_2_addbus_[6])
);
conv2d #("weight/conv2d_5/2_7.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_2_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_2_addbus_[7])
);
conv2d #("weight/conv2d_5/2_8.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_2_8(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[8]),
	.d_out(_2_addbus_[8])
);
conv2d #("weight/conv2d_5/2_9.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_2_9(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[9]),
	.d_out(_2_addbus_[9])
);
conv2d #("weight/conv2d_5/2_10.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_2_10(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[10]),
	.d_out(_2_addbus_[10])
);
conv2d #("weight/conv2d_5/2_11.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_2_11(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[11]),
	.d_out(_2_addbus_[11])
);
conv2d #("weight/conv2d_5/2_12.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_2_12(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[12]),
	.d_out(_2_addbus_[12])
);
conv2d #("weight/conv2d_5/2_13.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_2_13(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[13]),
	.d_out(_2_addbus_[13])
);
conv2d #("weight/conv2d_5/2_14.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_2_14(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[14]),
	.d_out(_2_addbus_[14])
);
conv2d #("weight/conv2d_5/2_15.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_2_15(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[15]),
	.d_out(_2_addbus_[15])
);
sum_16 #(3) sum_2( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[2]), 
        .data_in_0(_2_addbus_[0]), 
        .data_in_1(_2_addbus_[1]), 
        .data_in_2(_2_addbus_[2]), 
        .data_in_3(_2_addbus_[3]), 
        .data_in_4(_2_addbus_[4]), 
        .data_in_5(_2_addbus_[5]), 
        .data_in_6(_2_addbus_[6]), 
        .data_in_7(_2_addbus_[7]), 
        .data_in_8(_2_addbus_[8]), 
        .data_in_9(_2_addbus_[9]), 
        .data_in_10(_2_addbus_[10]), 
        .data_in_11(_2_addbus_[11]), 
        .data_in_12(_2_addbus_[12]), 
        .data_in_13(_2_addbus_[13]), 
        .data_in_14(_2_addbus_[14]), 
        .data_in_15(_2_addbus_[15]) 
); 
wire [31:0] _3_addbus_[15:0];    
conv2d #("weight/conv2d_5/3_0.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_3_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_3_addbus_[0])
);
conv2d #("weight/conv2d_5/3_1.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_3_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_3_addbus_[1])
);
conv2d #("weight/conv2d_5/3_2.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_3_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_3_addbus_[2])
);
conv2d #("weight/conv2d_5/3_3.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_3_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_3_addbus_[3])
);
conv2d #("weight/conv2d_5/3_4.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_3_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_3_addbus_[4])
);
conv2d #("weight/conv2d_5/3_5.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_3_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_3_addbus_[5])
);
conv2d #("weight/conv2d_5/3_6.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_3_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_3_addbus_[6])
);
conv2d #("weight/conv2d_5/3_7.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_3_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_3_addbus_[7])
);
conv2d #("weight/conv2d_5/3_8.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_3_8(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[8]),
	.d_out(_3_addbus_[8])
);
conv2d #("weight/conv2d_5/3_9.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_3_9(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[9]),
	.d_out(_3_addbus_[9])
);
conv2d #("weight/conv2d_5/3_10.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_3_10(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[10]),
	.d_out(_3_addbus_[10])
);
conv2d #("weight/conv2d_5/3_11.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_3_11(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[11]),
	.d_out(_3_addbus_[11])
);
conv2d #("weight/conv2d_5/3_12.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_3_12(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[12]),
	.d_out(_3_addbus_[12])
);
conv2d #("weight/conv2d_5/3_13.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_3_13(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[13]),
	.d_out(_3_addbus_[13])
);
conv2d #("weight/conv2d_5/3_14.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_3_14(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[14]),
	.d_out(_3_addbus_[14])
);
conv2d #("weight/conv2d_5/3_15.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_3_15(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[15]),
	.d_out(_3_addbus_[15])
);
sum_16 #(3) sum_3( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[3]), 
        .data_in_0(_3_addbus_[0]), 
        .data_in_1(_3_addbus_[1]), 
        .data_in_2(_3_addbus_[2]), 
        .data_in_3(_3_addbus_[3]), 
        .data_in_4(_3_addbus_[4]), 
        .data_in_5(_3_addbus_[5]), 
        .data_in_6(_3_addbus_[6]), 
        .data_in_7(_3_addbus_[7]), 
        .data_in_8(_3_addbus_[8]), 
        .data_in_9(_3_addbus_[9]), 
        .data_in_10(_3_addbus_[10]), 
        .data_in_11(_3_addbus_[11]), 
        .data_in_12(_3_addbus_[12]), 
        .data_in_13(_3_addbus_[13]), 
        .data_in_14(_3_addbus_[14]), 
        .data_in_15(_3_addbus_[15]) 
); 
wire [31:0] _4_addbus_[15:0];    
conv2d #("weight/conv2d_5/4_0.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_4_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_4_addbus_[0])
);
conv2d #("weight/conv2d_5/4_1.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_4_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_4_addbus_[1])
);
conv2d #("weight/conv2d_5/4_2.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_4_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_4_addbus_[2])
);
conv2d #("weight/conv2d_5/4_3.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_4_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_4_addbus_[3])
);
conv2d #("weight/conv2d_5/4_4.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_4_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_4_addbus_[4])
);
conv2d #("weight/conv2d_5/4_5.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_4_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_4_addbus_[5])
);
conv2d #("weight/conv2d_5/4_6.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_4_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_4_addbus_[6])
);
conv2d #("weight/conv2d_5/4_7.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_4_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_4_addbus_[7])
);
conv2d #("weight/conv2d_5/4_8.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_4_8(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[8]),
	.d_out(_4_addbus_[8])
);
conv2d #("weight/conv2d_5/4_9.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_4_9(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[9]),
	.d_out(_4_addbus_[9])
);
conv2d #("weight/conv2d_5/4_10.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_4_10(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[10]),
	.d_out(_4_addbus_[10])
);
conv2d #("weight/conv2d_5/4_11.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_4_11(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[11]),
	.d_out(_4_addbus_[11])
);
conv2d #("weight/conv2d_5/4_12.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_4_12(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[12]),
	.d_out(_4_addbus_[12])
);
conv2d #("weight/conv2d_5/4_13.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_4_13(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[13]),
	.d_out(_4_addbus_[13])
);
conv2d #("weight/conv2d_5/4_14.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_4_14(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[14]),
	.d_out(_4_addbus_[14])
);
conv2d #("weight/conv2d_5/4_15.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_4_15(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[15]),
	.d_out(_4_addbus_[15])
);
sum_16 #(3) sum_4( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[4]), 
        .data_in_0(_4_addbus_[0]), 
        .data_in_1(_4_addbus_[1]), 
        .data_in_2(_4_addbus_[2]), 
        .data_in_3(_4_addbus_[3]), 
        .data_in_4(_4_addbus_[4]), 
        .data_in_5(_4_addbus_[5]), 
        .data_in_6(_4_addbus_[6]), 
        .data_in_7(_4_addbus_[7]), 
        .data_in_8(_4_addbus_[8]), 
        .data_in_9(_4_addbus_[9]), 
        .data_in_10(_4_addbus_[10]), 
        .data_in_11(_4_addbus_[11]), 
        .data_in_12(_4_addbus_[12]), 
        .data_in_13(_4_addbus_[13]), 
        .data_in_14(_4_addbus_[14]), 
        .data_in_15(_4_addbus_[15]) 
); 
wire [31:0] _5_addbus_[15:0];    
conv2d #("weight/conv2d_5/5_0.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_5_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_5_addbus_[0])
);
conv2d #("weight/conv2d_5/5_1.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_5_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_5_addbus_[1])
);
conv2d #("weight/conv2d_5/5_2.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_5_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_5_addbus_[2])
);
conv2d #("weight/conv2d_5/5_3.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_5_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_5_addbus_[3])
);
conv2d #("weight/conv2d_5/5_4.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_5_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_5_addbus_[4])
);
conv2d #("weight/conv2d_5/5_5.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_5_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_5_addbus_[5])
);
conv2d #("weight/conv2d_5/5_6.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_5_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_5_addbus_[6])
);
conv2d #("weight/conv2d_5/5_7.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_5_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_5_addbus_[7])
);
conv2d #("weight/conv2d_5/5_8.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_5_8(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[8]),
	.d_out(_5_addbus_[8])
);
conv2d #("weight/conv2d_5/5_9.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_5_9(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[9]),
	.d_out(_5_addbus_[9])
);
conv2d #("weight/conv2d_5/5_10.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_5_10(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[10]),
	.d_out(_5_addbus_[10])
);
conv2d #("weight/conv2d_5/5_11.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_5_11(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[11]),
	.d_out(_5_addbus_[11])
);
conv2d #("weight/conv2d_5/5_12.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_5_12(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[12]),
	.d_out(_5_addbus_[12])
);
conv2d #("weight/conv2d_5/5_13.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_5_13(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[13]),
	.d_out(_5_addbus_[13])
);
conv2d #("weight/conv2d_5/5_14.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_5_14(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[14]),
	.d_out(_5_addbus_[14])
);
conv2d #("weight/conv2d_5/5_15.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_5_15(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[15]),
	.d_out(_5_addbus_[15])
);
sum_16 #(3) sum_5( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[5]), 
        .data_in_0(_5_addbus_[0]), 
        .data_in_1(_5_addbus_[1]), 
        .data_in_2(_5_addbus_[2]), 
        .data_in_3(_5_addbus_[3]), 
        .data_in_4(_5_addbus_[4]), 
        .data_in_5(_5_addbus_[5]), 
        .data_in_6(_5_addbus_[6]), 
        .data_in_7(_5_addbus_[7]), 
        .data_in_8(_5_addbus_[8]), 
        .data_in_9(_5_addbus_[9]), 
        .data_in_10(_5_addbus_[10]), 
        .data_in_11(_5_addbus_[11]), 
        .data_in_12(_5_addbus_[12]), 
        .data_in_13(_5_addbus_[13]), 
        .data_in_14(_5_addbus_[14]), 
        .data_in_15(_5_addbus_[15]) 
); 
wire [31:0] _6_addbus_[15:0];    
conv2d #("weight/conv2d_5/6_0.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_6_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_6_addbus_[0])
);
conv2d #("weight/conv2d_5/6_1.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_6_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_6_addbus_[1])
);
conv2d #("weight/conv2d_5/6_2.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_6_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_6_addbus_[2])
);
conv2d #("weight/conv2d_5/6_3.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_6_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_6_addbus_[3])
);
conv2d #("weight/conv2d_5/6_4.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_6_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_6_addbus_[4])
);
conv2d #("weight/conv2d_5/6_5.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_6_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_6_addbus_[5])
);
conv2d #("weight/conv2d_5/6_6.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_6_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_6_addbus_[6])
);
conv2d #("weight/conv2d_5/6_7.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_6_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_6_addbus_[7])
);
conv2d #("weight/conv2d_5/6_8.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_6_8(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[8]),
	.d_out(_6_addbus_[8])
);
conv2d #("weight/conv2d_5/6_9.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_6_9(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[9]),
	.d_out(_6_addbus_[9])
);
conv2d #("weight/conv2d_5/6_10.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_6_10(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[10]),
	.d_out(_6_addbus_[10])
);
conv2d #("weight/conv2d_5/6_11.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_6_11(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[11]),
	.d_out(_6_addbus_[11])
);
conv2d #("weight/conv2d_5/6_12.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_6_12(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[12]),
	.d_out(_6_addbus_[12])
);
conv2d #("weight/conv2d_5/6_13.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_6_13(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[13]),
	.d_out(_6_addbus_[13])
);
conv2d #("weight/conv2d_5/6_14.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_6_14(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[14]),
	.d_out(_6_addbus_[14])
);
conv2d #("weight/conv2d_5/6_15.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_6_15(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[15]),
	.d_out(_6_addbus_[15])
);
sum_16 #(3) sum_6( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[6]), 
        .data_in_0(_6_addbus_[0]), 
        .data_in_1(_6_addbus_[1]), 
        .data_in_2(_6_addbus_[2]), 
        .data_in_3(_6_addbus_[3]), 
        .data_in_4(_6_addbus_[4]), 
        .data_in_5(_6_addbus_[5]), 
        .data_in_6(_6_addbus_[6]), 
        .data_in_7(_6_addbus_[7]), 
        .data_in_8(_6_addbus_[8]), 
        .data_in_9(_6_addbus_[9]), 
        .data_in_10(_6_addbus_[10]), 
        .data_in_11(_6_addbus_[11]), 
        .data_in_12(_6_addbus_[12]), 
        .data_in_13(_6_addbus_[13]), 
        .data_in_14(_6_addbus_[14]), 
        .data_in_15(_6_addbus_[15]) 
); 
wire [31:0] _7_addbus_[15:0];    
conv2d #("weight/conv2d_5/7_0.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_7_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_7_addbus_[0])
);
conv2d #("weight/conv2d_5/7_1.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_7_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_7_addbus_[1])
);
conv2d #("weight/conv2d_5/7_2.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_7_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_7_addbus_[2])
);
conv2d #("weight/conv2d_5/7_3.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_7_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_7_addbus_[3])
);
conv2d #("weight/conv2d_5/7_4.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_7_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_7_addbus_[4])
);
conv2d #("weight/conv2d_5/7_5.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_7_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_7_addbus_[5])
);
conv2d #("weight/conv2d_5/7_6.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_7_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_7_addbus_[6])
);
conv2d #("weight/conv2d_5/7_7.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_7_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_7_addbus_[7])
);
conv2d #("weight/conv2d_5/7_8.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_7_8(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[8]),
	.d_out(_7_addbus_[8])
);
conv2d #("weight/conv2d_5/7_9.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_7_9(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[9]),
	.d_out(_7_addbus_[9])
);
conv2d #("weight/conv2d_5/7_10.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_7_10(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[10]),
	.d_out(_7_addbus_[10])
);
conv2d #("weight/conv2d_5/7_11.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_7_11(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[11]),
	.d_out(_7_addbus_[11])
);
conv2d #("weight/conv2d_5/7_12.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_7_12(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[12]),
	.d_out(_7_addbus_[12])
);
conv2d #("weight/conv2d_5/7_13.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_7_13(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[13]),
	.d_out(_7_addbus_[13])
);
conv2d #("weight/conv2d_5/7_14.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_7_14(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[14]),
	.d_out(_7_addbus_[14])
);
conv2d #("weight/conv2d_5/7_15.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_7_15(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[15]),
	.d_out(_7_addbus_[15])
);
sum_16 #(3) sum_7( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[7]), 
        .data_in_0(_7_addbus_[0]), 
        .data_in_1(_7_addbus_[1]), 
        .data_in_2(_7_addbus_[2]), 
        .data_in_3(_7_addbus_[3]), 
        .data_in_4(_7_addbus_[4]), 
        .data_in_5(_7_addbus_[5]), 
        .data_in_6(_7_addbus_[6]), 
        .data_in_7(_7_addbus_[7]), 
        .data_in_8(_7_addbus_[8]), 
        .data_in_9(_7_addbus_[9]), 
        .data_in_10(_7_addbus_[10]), 
        .data_in_11(_7_addbus_[11]), 
        .data_in_12(_7_addbus_[12]), 
        .data_in_13(_7_addbus_[13]), 
        .data_in_14(_7_addbus_[14]), 
        .data_in_15(_7_addbus_[15]) 
); 
wire [31:0] _8_addbus_[15:0];    
conv2d #("weight/conv2d_5/8_0.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_8_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_8_addbus_[0])
);
conv2d #("weight/conv2d_5/8_1.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_8_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_8_addbus_[1])
);
conv2d #("weight/conv2d_5/8_2.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_8_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_8_addbus_[2])
);
conv2d #("weight/conv2d_5/8_3.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_8_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_8_addbus_[3])
);
conv2d #("weight/conv2d_5/8_4.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_8_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_8_addbus_[4])
);
conv2d #("weight/conv2d_5/8_5.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_8_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_8_addbus_[5])
);
conv2d #("weight/conv2d_5/8_6.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_8_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_8_addbus_[6])
);
conv2d #("weight/conv2d_5/8_7.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_8_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_8_addbus_[7])
);
conv2d #("weight/conv2d_5/8_8.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_8_8(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[8]),
	.d_out(_8_addbus_[8])
);
conv2d #("weight/conv2d_5/8_9.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_8_9(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[9]),
	.d_out(_8_addbus_[9])
);
conv2d #("weight/conv2d_5/8_10.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_8_10(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[10]),
	.d_out(_8_addbus_[10])
);
conv2d #("weight/conv2d_5/8_11.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_8_11(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[11]),
	.d_out(_8_addbus_[11])
);
conv2d #("weight/conv2d_5/8_12.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_8_12(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[12]),
	.d_out(_8_addbus_[12])
);
conv2d #("weight/conv2d_5/8_13.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_8_13(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[13]),
	.d_out(_8_addbus_[13])
);
conv2d #("weight/conv2d_5/8_14.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_8_14(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[14]),
	.d_out(_8_addbus_[14])
);
conv2d #("weight/conv2d_5/8_15.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_8_15(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[15]),
	.d_out(_8_addbus_[15])
);
sum_16 #(3) sum_8( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[8]), 
        .data_in_0(_8_addbus_[0]), 
        .data_in_1(_8_addbus_[1]), 
        .data_in_2(_8_addbus_[2]), 
        .data_in_3(_8_addbus_[3]), 
        .data_in_4(_8_addbus_[4]), 
        .data_in_5(_8_addbus_[5]), 
        .data_in_6(_8_addbus_[6]), 
        .data_in_7(_8_addbus_[7]), 
        .data_in_8(_8_addbus_[8]), 
        .data_in_9(_8_addbus_[9]), 
        .data_in_10(_8_addbus_[10]), 
        .data_in_11(_8_addbus_[11]), 
        .data_in_12(_8_addbus_[12]), 
        .data_in_13(_8_addbus_[13]), 
        .data_in_14(_8_addbus_[14]), 
        .data_in_15(_8_addbus_[15]) 
); 
wire [31:0] _9_addbus_[15:0];    
conv2d #("weight/conv2d_5/9_0.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_9_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_9_addbus_[0])
);
conv2d #("weight/conv2d_5/9_1.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_9_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_9_addbus_[1])
);
conv2d #("weight/conv2d_5/9_2.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_9_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_9_addbus_[2])
);
conv2d #("weight/conv2d_5/9_3.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_9_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_9_addbus_[3])
);
conv2d #("weight/conv2d_5/9_4.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_9_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_9_addbus_[4])
);
conv2d #("weight/conv2d_5/9_5.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_9_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_9_addbus_[5])
);
conv2d #("weight/conv2d_5/9_6.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_9_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_9_addbus_[6])
);
conv2d #("weight/conv2d_5/9_7.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_9_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_9_addbus_[7])
);
conv2d #("weight/conv2d_5/9_8.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_9_8(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[8]),
	.d_out(_9_addbus_[8])
);
conv2d #("weight/conv2d_5/9_9.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_9_9(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[9]),
	.d_out(_9_addbus_[9])
);
conv2d #("weight/conv2d_5/9_10.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_9_10(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[10]),
	.d_out(_9_addbus_[10])
);
conv2d #("weight/conv2d_5/9_11.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_9_11(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[11]),
	.d_out(_9_addbus_[11])
);
conv2d #("weight/conv2d_5/9_12.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_9_12(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[12]),
	.d_out(_9_addbus_[12])
);
conv2d #("weight/conv2d_5/9_13.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_9_13(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[13]),
	.d_out(_9_addbus_[13])
);
conv2d #("weight/conv2d_5/9_14.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_9_14(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[14]),
	.d_out(_9_addbus_[14])
);
conv2d #("weight/conv2d_5/9_15.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_9_15(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[15]),
	.d_out(_9_addbus_[15])
);
sum_16 #(3) sum_9( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[9]), 
        .data_in_0(_9_addbus_[0]), 
        .data_in_1(_9_addbus_[1]), 
        .data_in_2(_9_addbus_[2]), 
        .data_in_3(_9_addbus_[3]), 
        .data_in_4(_9_addbus_[4]), 
        .data_in_5(_9_addbus_[5]), 
        .data_in_6(_9_addbus_[6]), 
        .data_in_7(_9_addbus_[7]), 
        .data_in_8(_9_addbus_[8]), 
        .data_in_9(_9_addbus_[9]), 
        .data_in_10(_9_addbus_[10]), 
        .data_in_11(_9_addbus_[11]), 
        .data_in_12(_9_addbus_[12]), 
        .data_in_13(_9_addbus_[13]), 
        .data_in_14(_9_addbus_[14]), 
        .data_in_15(_9_addbus_[15]) 
); 
wire [31:0] _10_addbus_[15:0];    
conv2d #("weight/conv2d_5/10_0.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_10_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_10_addbus_[0])
);
conv2d #("weight/conv2d_5/10_1.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_10_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_10_addbus_[1])
);
conv2d #("weight/conv2d_5/10_2.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_10_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_10_addbus_[2])
);
conv2d #("weight/conv2d_5/10_3.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_10_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_10_addbus_[3])
);
conv2d #("weight/conv2d_5/10_4.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_10_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_10_addbus_[4])
);
conv2d #("weight/conv2d_5/10_5.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_10_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_10_addbus_[5])
);
conv2d #("weight/conv2d_5/10_6.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_10_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_10_addbus_[6])
);
conv2d #("weight/conv2d_5/10_7.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_10_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_10_addbus_[7])
);
conv2d #("weight/conv2d_5/10_8.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_10_8(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[8]),
	.d_out(_10_addbus_[8])
);
conv2d #("weight/conv2d_5/10_9.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_10_9(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[9]),
	.d_out(_10_addbus_[9])
);
conv2d #("weight/conv2d_5/10_10.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_10_10(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[10]),
	.d_out(_10_addbus_[10])
);
conv2d #("weight/conv2d_5/10_11.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_10_11(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[11]),
	.d_out(_10_addbus_[11])
);
conv2d #("weight/conv2d_5/10_12.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_10_12(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[12]),
	.d_out(_10_addbus_[12])
);
conv2d #("weight/conv2d_5/10_13.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_10_13(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[13]),
	.d_out(_10_addbus_[13])
);
conv2d #("weight/conv2d_5/10_14.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_10_14(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[14]),
	.d_out(_10_addbus_[14])
);
conv2d #("weight/conv2d_5/10_15.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_10_15(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[15]),
	.d_out(_10_addbus_[15])
);
sum_16 #(3) sum_10( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[10]), 
        .data_in_0(_10_addbus_[0]), 
        .data_in_1(_10_addbus_[1]), 
        .data_in_2(_10_addbus_[2]), 
        .data_in_3(_10_addbus_[3]), 
        .data_in_4(_10_addbus_[4]), 
        .data_in_5(_10_addbus_[5]), 
        .data_in_6(_10_addbus_[6]), 
        .data_in_7(_10_addbus_[7]), 
        .data_in_8(_10_addbus_[8]), 
        .data_in_9(_10_addbus_[9]), 
        .data_in_10(_10_addbus_[10]), 
        .data_in_11(_10_addbus_[11]), 
        .data_in_12(_10_addbus_[12]), 
        .data_in_13(_10_addbus_[13]), 
        .data_in_14(_10_addbus_[14]), 
        .data_in_15(_10_addbus_[15]) 
); 
wire [31:0] _11_addbus_[15:0];    
conv2d #("weight/conv2d_5/11_0.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_11_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_11_addbus_[0])
);
conv2d #("weight/conv2d_5/11_1.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_11_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_11_addbus_[1])
);
conv2d #("weight/conv2d_5/11_2.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_11_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_11_addbus_[2])
);
conv2d #("weight/conv2d_5/11_3.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_11_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_11_addbus_[3])
);
conv2d #("weight/conv2d_5/11_4.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_11_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_11_addbus_[4])
);
conv2d #("weight/conv2d_5/11_5.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_11_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_11_addbus_[5])
);
conv2d #("weight/conv2d_5/11_6.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_11_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_11_addbus_[6])
);
conv2d #("weight/conv2d_5/11_7.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_11_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_11_addbus_[7])
);
conv2d #("weight/conv2d_5/11_8.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_11_8(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[8]),
	.d_out(_11_addbus_[8])
);
conv2d #("weight/conv2d_5/11_9.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_11_9(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[9]),
	.d_out(_11_addbus_[9])
);
conv2d #("weight/conv2d_5/11_10.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_11_10(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[10]),
	.d_out(_11_addbus_[10])
);
conv2d #("weight/conv2d_5/11_11.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_11_11(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[11]),
	.d_out(_11_addbus_[11])
);
conv2d #("weight/conv2d_5/11_12.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_11_12(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[12]),
	.d_out(_11_addbus_[12])
);
conv2d #("weight/conv2d_5/11_13.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_11_13(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[13]),
	.d_out(_11_addbus_[13])
);
conv2d #("weight/conv2d_5/11_14.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_11_14(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[14]),
	.d_out(_11_addbus_[14])
);
conv2d #("weight/conv2d_5/11_15.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_11_15(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[15]),
	.d_out(_11_addbus_[15])
);
sum_16 #(3) sum_11( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[11]), 
        .data_in_0(_11_addbus_[0]), 
        .data_in_1(_11_addbus_[1]), 
        .data_in_2(_11_addbus_[2]), 
        .data_in_3(_11_addbus_[3]), 
        .data_in_4(_11_addbus_[4]), 
        .data_in_5(_11_addbus_[5]), 
        .data_in_6(_11_addbus_[6]), 
        .data_in_7(_11_addbus_[7]), 
        .data_in_8(_11_addbus_[8]), 
        .data_in_9(_11_addbus_[9]), 
        .data_in_10(_11_addbus_[10]), 
        .data_in_11(_11_addbus_[11]), 
        .data_in_12(_11_addbus_[12]), 
        .data_in_13(_11_addbus_[13]), 
        .data_in_14(_11_addbus_[14]), 
        .data_in_15(_11_addbus_[15]) 
); 
wire [31:0] _12_addbus_[15:0];    
conv2d #("weight/conv2d_5/12_0.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_12_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_12_addbus_[0])
);
conv2d #("weight/conv2d_5/12_1.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_12_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_12_addbus_[1])
);
conv2d #("weight/conv2d_5/12_2.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_12_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_12_addbus_[2])
);
conv2d #("weight/conv2d_5/12_3.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_12_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_12_addbus_[3])
);
conv2d #("weight/conv2d_5/12_4.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_12_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_12_addbus_[4])
);
conv2d #("weight/conv2d_5/12_5.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_12_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_12_addbus_[5])
);
conv2d #("weight/conv2d_5/12_6.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_12_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_12_addbus_[6])
);
conv2d #("weight/conv2d_5/12_7.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_12_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_12_addbus_[7])
);
conv2d #("weight/conv2d_5/12_8.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_12_8(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[8]),
	.d_out(_12_addbus_[8])
);
conv2d #("weight/conv2d_5/12_9.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_12_9(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[9]),
	.d_out(_12_addbus_[9])
);
conv2d #("weight/conv2d_5/12_10.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_12_10(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[10]),
	.d_out(_12_addbus_[10])
);
conv2d #("weight/conv2d_5/12_11.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_12_11(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[11]),
	.d_out(_12_addbus_[11])
);
conv2d #("weight/conv2d_5/12_12.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_12_12(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[12]),
	.d_out(_12_addbus_[12])
);
conv2d #("weight/conv2d_5/12_13.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_12_13(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[13]),
	.d_out(_12_addbus_[13])
);
conv2d #("weight/conv2d_5/12_14.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_12_14(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[14]),
	.d_out(_12_addbus_[14])
);
conv2d #("weight/conv2d_5/12_15.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_12_15(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[15]),
	.d_out(_12_addbus_[15])
);
sum_16 #(3) sum_12( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[12]), 
        .data_in_0(_12_addbus_[0]), 
        .data_in_1(_12_addbus_[1]), 
        .data_in_2(_12_addbus_[2]), 
        .data_in_3(_12_addbus_[3]), 
        .data_in_4(_12_addbus_[4]), 
        .data_in_5(_12_addbus_[5]), 
        .data_in_6(_12_addbus_[6]), 
        .data_in_7(_12_addbus_[7]), 
        .data_in_8(_12_addbus_[8]), 
        .data_in_9(_12_addbus_[9]), 
        .data_in_10(_12_addbus_[10]), 
        .data_in_11(_12_addbus_[11]), 
        .data_in_12(_12_addbus_[12]), 
        .data_in_13(_12_addbus_[13]), 
        .data_in_14(_12_addbus_[14]), 
        .data_in_15(_12_addbus_[15]) 
); 
wire [31:0] _13_addbus_[15:0];    
conv2d #("weight/conv2d_5/13_0.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_13_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_13_addbus_[0])
);
conv2d #("weight/conv2d_5/13_1.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_13_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_13_addbus_[1])
);
conv2d #("weight/conv2d_5/13_2.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_13_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_13_addbus_[2])
);
conv2d #("weight/conv2d_5/13_3.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_13_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_13_addbus_[3])
);
conv2d #("weight/conv2d_5/13_4.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_13_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_13_addbus_[4])
);
conv2d #("weight/conv2d_5/13_5.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_13_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_13_addbus_[5])
);
conv2d #("weight/conv2d_5/13_6.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_13_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_13_addbus_[6])
);
conv2d #("weight/conv2d_5/13_7.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_13_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_13_addbus_[7])
);
conv2d #("weight/conv2d_5/13_8.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_13_8(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[8]),
	.d_out(_13_addbus_[8])
);
conv2d #("weight/conv2d_5/13_9.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_13_9(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[9]),
	.d_out(_13_addbus_[9])
);
conv2d #("weight/conv2d_5/13_10.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_13_10(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[10]),
	.d_out(_13_addbus_[10])
);
conv2d #("weight/conv2d_5/13_11.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_13_11(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[11]),
	.d_out(_13_addbus_[11])
);
conv2d #("weight/conv2d_5/13_12.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_13_12(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[12]),
	.d_out(_13_addbus_[12])
);
conv2d #("weight/conv2d_5/13_13.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_13_13(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[13]),
	.d_out(_13_addbus_[13])
);
conv2d #("weight/conv2d_5/13_14.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_13_14(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[14]),
	.d_out(_13_addbus_[14])
);
conv2d #("weight/conv2d_5/13_15.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_13_15(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[15]),
	.d_out(_13_addbus_[15])
);
sum_16 #(3) sum_13( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[13]), 
        .data_in_0(_13_addbus_[0]), 
        .data_in_1(_13_addbus_[1]), 
        .data_in_2(_13_addbus_[2]), 
        .data_in_3(_13_addbus_[3]), 
        .data_in_4(_13_addbus_[4]), 
        .data_in_5(_13_addbus_[5]), 
        .data_in_6(_13_addbus_[6]), 
        .data_in_7(_13_addbus_[7]), 
        .data_in_8(_13_addbus_[8]), 
        .data_in_9(_13_addbus_[9]), 
        .data_in_10(_13_addbus_[10]), 
        .data_in_11(_13_addbus_[11]), 
        .data_in_12(_13_addbus_[12]), 
        .data_in_13(_13_addbus_[13]), 
        .data_in_14(_13_addbus_[14]), 
        .data_in_15(_13_addbus_[15]) 
); 
wire [31:0] _14_addbus_[15:0];    
conv2d #("weight/conv2d_5/14_0.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_14_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_14_addbus_[0])
);
conv2d #("weight/conv2d_5/14_1.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_14_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_14_addbus_[1])
);
conv2d #("weight/conv2d_5/14_2.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_14_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_14_addbus_[2])
);
conv2d #("weight/conv2d_5/14_3.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_14_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_14_addbus_[3])
);
conv2d #("weight/conv2d_5/14_4.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_14_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_14_addbus_[4])
);
conv2d #("weight/conv2d_5/14_5.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_14_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_14_addbus_[5])
);
conv2d #("weight/conv2d_5/14_6.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_14_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_14_addbus_[6])
);
conv2d #("weight/conv2d_5/14_7.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_14_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_14_addbus_[7])
);
conv2d #("weight/conv2d_5/14_8.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_14_8(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[8]),
	.d_out(_14_addbus_[8])
);
conv2d #("weight/conv2d_5/14_9.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_14_9(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[9]),
	.d_out(_14_addbus_[9])
);
conv2d #("weight/conv2d_5/14_10.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_14_10(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[10]),
	.d_out(_14_addbus_[10])
);
conv2d #("weight/conv2d_5/14_11.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_14_11(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[11]),
	.d_out(_14_addbus_[11])
);
conv2d #("weight/conv2d_5/14_12.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_14_12(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[12]),
	.d_out(_14_addbus_[12])
);
conv2d #("weight/conv2d_5/14_13.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_14_13(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[13]),
	.d_out(_14_addbus_[13])
);
conv2d #("weight/conv2d_5/14_14.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_14_14(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[14]),
	.d_out(_14_addbus_[14])
);
conv2d #("weight/conv2d_5/14_15.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_14_15(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[15]),
	.d_out(_14_addbus_[15])
);
sum_16 #(3) sum_14( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[14]), 
        .data_in_0(_14_addbus_[0]), 
        .data_in_1(_14_addbus_[1]), 
        .data_in_2(_14_addbus_[2]), 
        .data_in_3(_14_addbus_[3]), 
        .data_in_4(_14_addbus_[4]), 
        .data_in_5(_14_addbus_[5]), 
        .data_in_6(_14_addbus_[6]), 
        .data_in_7(_14_addbus_[7]), 
        .data_in_8(_14_addbus_[8]), 
        .data_in_9(_14_addbus_[9]), 
        .data_in_10(_14_addbus_[10]), 
        .data_in_11(_14_addbus_[11]), 
        .data_in_12(_14_addbus_[12]), 
        .data_in_13(_14_addbus_[13]), 
        .data_in_14(_14_addbus_[14]), 
        .data_in_15(_14_addbus_[15]) 
); 
wire [31:0] _15_addbus_[15:0];    
conv2d #("weight/conv2d_5/15_0.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_15_0(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[0]),
	.d_out(_15_addbus_[0])
);
conv2d #("weight/conv2d_5/15_1.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_15_1(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[1]),
	.d_out(_15_addbus_[1])
);
conv2d #("weight/conv2d_5/15_2.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_15_2(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[2]),
	.d_out(_15_addbus_[2])
);
conv2d #("weight/conv2d_5/15_3.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_15_3(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[3]),
	.d_out(_15_addbus_[3])
);
conv2d #("weight/conv2d_5/15_4.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_15_4(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[4]),
	.d_out(_15_addbus_[4])
);
conv2d #("weight/conv2d_5/15_5.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_15_5(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[5]),
	.d_out(_15_addbus_[5])
);
conv2d #("weight/conv2d_5/15_6.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_15_6(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[6]),
	.d_out(_15_addbus_[6])
);
conv2d #("weight/conv2d_5/15_7.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_15_7(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[7]),
	.d_out(_15_addbus_[7])
);
conv2d #("weight/conv2d_5/15_8.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_15_8(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[8]),
	.d_out(_15_addbus_[8])
);
conv2d #("weight/conv2d_5/15_9.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_15_9(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[9]),
	.d_out(_15_addbus_[9])
);
conv2d #("weight/conv2d_5/15_10.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_15_10(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[10]),
	.d_out(_15_addbus_[10])
);
conv2d #("weight/conv2d_5/15_11.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_15_11(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[11]),
	.d_out(_15_addbus_[11])
);
conv2d #("weight/conv2d_5/15_12.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_15_12(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[12]),
	.d_out(_15_addbus_[12])
);
conv2d #("weight/conv2d_5/15_13.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_15_13(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[13]),
	.d_out(_15_addbus_[13])
);
conv2d #("weight/conv2d_5/15_14.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_15_14(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[14]),
	.d_out(_15_addbus_[14])
);
conv2d #("weight/conv2d_5/15_15.txt", 0 /*dont use relu*/, 1, 1, 3, 3) conv2d_15_15(
	.clk(clk),
	.rst(rst),
	.input_valid(input_valid),
	.load(load),
	.load_success(),
	.output_valid(),
	.sof(sof),
	.o_sof(),
	.d_in(d_in[15]),
	.d_out(_15_addbus_[15])
);
sum_16 #(3) sum_15( 
        .clk(clk), 
        .rst(rst), 
        .input_valid(output_valid_affter_conv), 
        .data_out(d_out[15]), 
        .data_in_0(_15_addbus_[0]), 
        .data_in_1(_15_addbus_[1]), 
        .data_in_2(_15_addbus_[2]), 
        .data_in_3(_15_addbus_[3]), 
        .data_in_4(_15_addbus_[4]), 
        .data_in_5(_15_addbus_[5]), 
        .data_in_6(_15_addbus_[6]), 
        .data_in_7(_15_addbus_[7]), 
        .data_in_8(_15_addbus_[8]), 
        .data_in_9(_15_addbus_[9]), 
        .data_in_10(_15_addbus_[10]), 
        .data_in_11(_15_addbus_[11]), 
        .data_in_12(_15_addbus_[12]), 
        .data_in_13(_15_addbus_[13]), 
        .data_in_14(_15_addbus_[14]), 
        .data_in_15(_15_addbus_[15]) 
); 
endmodule